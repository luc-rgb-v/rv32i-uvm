`ifndef BUS_DEFINES
`define BUS_DEFINES

  `define NO_OF_TRANSACTIONS 1000
  `define BUS_ADDR_WIDTH 32
  `define BUS_DATA_WIDTH 32

`endif
